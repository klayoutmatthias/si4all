* Netlist after simplification

* cell RINGO
* pin FB
* pin VDD
* pin OUT
* pin ENABLE
* pin BULK,VSS
.SUBCKT RINGO FB VDD OUT ENABLE BULK|VSS
* cell instance $1 r0 *1 1.8,0
X$1 VDD \$1 BULK|VSS VDD FB ENABLE BULK|VSS ND2X1
* cell instance $2 r0 *1 4.2,0
X$2 VDD \$2 BULK|VSS VDD \$1 BULK|VSS INVX1
* cell instance $3 r0 *1 6,0
X$3 VDD \$3 BULK|VSS VDD \$2 BULK|VSS INVX1
* cell instance $4 r0 *1 7.8,0
X$4 VDD \$4 BULK|VSS VDD \$3 BULK|VSS INVX1
* cell instance $5 r0 *1 9.6,0
X$5 VDD \$5 BULK|VSS VDD \$4 BULK|VSS INVX1
* cell instance $6 r0 *1 11.4,0
X$6 VDD \$6 BULK|VSS VDD \$5 BULK|VSS INVX1
* cell instance $7 r0 *1 13.2,0
X$7 VDD \$7 BULK|VSS VDD \$6 BULK|VSS INVX1
* cell instance $8 r0 *1 15,0
X$8 VDD \$8 BULK|VSS VDD \$7 BULK|VSS INVX1
* cell instance $9 r0 *1 16.8,0
X$9 VDD \$9 BULK|VSS VDD \$8 BULK|VSS INVX1
* cell instance $10 r0 *1 18.6,0
X$10 VDD \$10 BULK|VSS VDD \$9 BULK|VSS INVX1
* cell instance $11 r0 *1 20.4,0
X$11 VDD FB BULK|VSS VDD \$10 BULK|VSS INVX1
* cell instance $12 r0 *1 22.2,0
X$12 VDD OUT BULK|VSS VDD FB BULK|VSS INVX1
.ENDS RINGO

* cell ND2X1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin B
* pin A
* pin BULK
.SUBCKT ND2X1 VDD OUT VSS \$4 B A BULK
* device instance $1 0.85,5.8 LVPMOS
M$1 OUT A VDD \$4 MLVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 1.55,5.8 LVPMOS
M$2 VDD B OUT \$4 MLVPMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 0.85,2.135 LVNMOS
M$3 VSS A \$I3 BULK MLVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U
+ PD=1.4U
* device instance $4 1.55,2.135 LVNMOS
M$4 \$I3 B OUT BULK MLVNMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U
+ PD=2.75U
.ENDS ND2X1

* cell INVX1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin IN
* pin BULK
.SUBCKT INVX1 VDD OUT VSS \$4 IN BULK
* device instance $1 0.85,5.8 LVPMOS
M$1 VDD IN OUT \$4 MLVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U
+ PD=3.85U
* device instance $2 0.85,2.135 LVNMOS
M$2 VSS IN OUT BULK MLVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
.ENDS INVX1
